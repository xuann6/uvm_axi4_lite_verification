
package axi4_lite_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // =========================================================================
    // Parameters
    // =========================================================================
    parameter int unsigned ADDR_WIDTH = 32;
    parameter int unsigned DATA_WIDTH = 32;
    parameter int unsigned STRB_WIDTH = DATA_WIDTH / 8;   // 4

    parameter int unsigned NUM_REGS  = 16;
    parameter int unsigned REG_BYTES = NUM_REGS * 4;      // 64 = 0x40
    parameter logic [ADDR_WIDTH-1:0] REG_BASE = 32'h0000_0000;
    parameter logic [ADDR_WIDTH-1:0] REG_HIGH = 32'h0000_003C;  // last valid addr

    parameter int unsigned CLK_PERIOD_NS    = 10;
    parameter int unsigned HANDSHAKE_TIMEOUT = 100;

    // =========================================================================
    // Enumerations
    // =========================================================================

    // Transaction type
    typedef enum logic {
        WRITE = 1'b0,
        READ  = 1'b1
    } trans_type_e;

    // AXI4-Lite response codes
    // IMPORTANT: SLVERR is 2'b10 per the AXI specification (Table A1-4).
    // This must match the DUT's RESP_SLVERR = 2'b10.
    typedef enum logic [1:0] {
        RESP_OKAY   = 2'b00,   // Normal successful completion
        RESP_EXOKAY = 2'b01,   // Exclusive OK (not generated by this slave)
        RESP_SLVERR = 2'b10,   // Slave error (out-of-range / unaligned address)
        RESP_DECERR = 2'b11    // Decode error (not generated by this slave)
    } axi_resp_e;

    // =========================================================================
    // Typedefs
    // =========================================================================
    typedef logic [ADDR_WIDTH-1:0] axi_addr_t;
    typedef logic [DATA_WIDTH-1:0] axi_data_t;
    typedef logic [STRB_WIDTH-1:0] axi_strb_t;
    typedef logic [1:0]            axi_resp_t;

    // =========================================================================
    // TB source file includes (strict bottom-up dependency order)
    // =========================================================================

    // Layer 1 – Transaction (no TB dependencies)
    `include "sequences/axi4_lite_transaction.sv"

    // Layer 2 – Sequences (depend on transaction)
    `include "sequences/axi4_lite_sequences.sv"

    // Layer 3 – Agent components (depend on transaction)
    `include "agents/axi4_lite_driver.sv"
    `include "agents/axi4_lite_monitor.sv"
    `include "agents/axi4_lite_scoreboard.sv"
    `include "agents/axi4_lite_coverage.sv"

    // Layer 4 – Agent (sequencer class also lives inside this file)
    `include "agents/axi4_lite_agent.sv"

    // Layer 5 – Environment
    `include "axi4_lite_env.sv"

    // Layer 6 – Tests
    `include "tests/axi4_lite_test.sv"

endpackage : axi4_lite_pkg
